library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Pipeline is

end Pipeline;

architecture behavior of Pipeline is
begin
end architecture behavior;
